module nor_gate(in1,in2,out);
  
  input in1,in2;
  output out;
  
  assign = in1 & in2;
endmodule

  
  
